module VexRiscvAxiLite (
    input aclk,
    input aresetn,

    output logic[ADDR_WIDTH-1:0]             i_m_axil_awaddr,
    output logic[2:0]                        i_m_axil_awprot,
    output logic                             i_m_axil_awvalid,
    input logic                              i_m_axil_awready,
    output logic[DATA_WIDTH-1:0]             i_m_axil_wdata,
    output logic[STRB_WIDTH-1:0]             i_m_axil_wstrb,
    output logic                             i_m_axil_wvalid,
    input logic                              i_m_axil_wready,
    input logic [1:0]                        i_m_axil_bresp,
    input logic                              i_m_axil_bvalid,
    output logic                             i_m_axil_bready,
    output logic[ADDR_WIDTH-1:0]             i_m_axil_araddr,
    output logic[2:0]                        i_m_axil_arprot,
    output logic                             i_m_axil_arvalid,
    input logic                              i_m_axil_arready,
    input logic [DATA_WIDTH-1:0]             i_m_axil_rdata,
    input logic [1:0]                        i_m_axil_rresp,
    input logic                              i_m_axil_rvalid,
    output logic                             i_m_axil_rready,

    output logic[ADDR_WIDTH-1:0]             d_m_axil_awaddr,
    output logic[2:0]                        d_m_axil_awprot,
    output logic                             d_m_axil_awvalid,
    input logic                              d_m_axil_awready,
    output logic[DATA_WIDTH-1:0]             d_m_axil_wdata,
    output logic[STRB_WIDTH-1:0]             d_m_axil_wstrb,
    output logic                             d_m_axil_wvalid,
    input logic                              d_m_axil_wready,
    input logic [1:0]                        d_m_axil_bresp,
    input logic                              d_m_axil_bvalid,
    output logic                             d_m_axil_bready,
    output logic[ADDR_WIDTH-1:0]             d_m_axil_araddr,
    output logic[2:0]                        d_m_axil_arprot,
    output logic                             d_m_axil_arvalid,
    input logic                              d_m_axil_arready,
    input logic [DATA_WIDTH-1:0]             d_m_axil_rdata,
    input logic [1:0]                        d_m_axil_rresp,
    input logic                              d_m_axil_rvalid,
    output logic                             d_m_axil_rready
);

axi_axil_adapter IAdapter 
(
    
);

VexRiscvAxi4 VexCPU 
(
    .timerInterrupt(?),
    .externalInterrupt(?),
    .softwareInterrupt(?),
    .debug_bus_cmd_valid(?),
    .debug_bus_cmd_ready(?),
    .debug_bus_cmd_payload_wr(?),
    .debug_bus_cmd_payload_address(?),
    .debug_bus_cmd_payload_data(?),
    .debug_bus_rsp_data(?),
    .debug_resetOut(?),
    
    .iBusAxi_ar_valid(),
    .iBusAxi_ar_ready(),
    .iBusAxi_ar_payload_addr(),
    .iBusAxi_ar_payload_id(),
    .iBusAxi_ar_payload_region(),
    .iBusAxi_ar_payload_len(),
    .iBusAxi_ar_payload_size(),
    .iBusAxi_ar_payload_burst(),
    .iBusAxi_ar_payload_lock(),
    .iBusAxi_ar_payload_cache(),
    .iBusAxi_ar_payload_qos(),
    .iBusAxi_ar_payload_prot(),
    .iBusAxi_r_valid(),
    .iBusAxi_r_ready(),
    .iBusAxi_r_payload_data(),
    .iBusAxi_r_payload_id(),
    .iBusAxi_r_payload_resp(),
    .iBusAxi_r_payload_last(),
    .dBusAxi_aw_valid(),
    .dBusAxi_aw_ready(),
    .dBusAxi_aw_payload_addr(),
    .dBusAxi_aw_payload_id(),
    .dBusAxi_aw_payload_region(),
    .dBusAxi_aw_payload_len(),
    .dBusAxi_aw_payload_size(),
    .dBusAxi_aw_payload_burst(),
    .dBusAxi_aw_payload_lock(),
    .dBusAxi_aw_payload_cache(),
    .dBusAxi_aw_payload_qos(),
    .dBusAxi_aw_payload_prot(),
    .dBusAxi_w_valid(),
    .dBusAxi_w_ready(),
    .dBusAxi_w_payload_data(),
    .dBusAxi_w_payload_strb(),
    .dBusAxi_w_payload_last(),
    .dBusAxi_b_valid(),
    .dBusAxi_b_ready(),
    .dBusAxi_b_payload_id(),
    .dBusAxi_b_payload_resp(),
    .dBusAxi_ar_valid(),
    .dBusAxi_ar_ready(),
    .dBusAxi_ar_payload_addr(),
    .dBusAxi_ar_payload_id(),
    .dBusAxi_ar_payload_region(),
    .dBusAxi_ar_payload_len(),
    .dBusAxi_ar_payload_size(),
    .dBusAxi_ar_payload_burst(),
    .dBusAxi_ar_payload_lock(),
    .dBusAxi_ar_payload_cache(),
    .dBusAxi_ar_payload_qos(),
    .dBusAxi_ar_payload_prot(),
    .dBusAxi_r_valid(),
    .dBusAxi_r_ready(),
    .dBusAxi_r_payload_data(),
    .dBusAxi_r_payload_id(),
    .dBusAxi_r_payload_resp(),
    .dBusAxi_r_payload_last(),
    .clk(),
    .reset(),
    .debugReset()
);
    
endmodule