module VexRiscvAxiLite (
    input aclk,
    input aresetn,

    output logic[ADDR_WIDTH-1:0]             i_m_axil_awaddr,
    output logic[2:0]                        i_m_axil_awprot,
    output logic                             i_m_axil_awvalid,
    input logic                              i_m_axil_awready,
    output logic[DATA_WIDTH-1:0]             i_m_axil_wdata,
    output logic[STRB_WIDTH-1:0]             i_m_axil_wstrb,
    output logic                             i_m_axil_wvalid,
    input logic                              i_m_axil_wready,
    input logic [1:0]                        i_m_axil_bresp,
    input logic                              i_m_axil_bvalid,
    output logic                             i_m_axil_bready,
    output logic[ADDR_WIDTH-1:0]             i_m_axil_araddr,
    output logic[2:0]                        i_m_axil_arprot,
    output logic                             i_m_axil_arvalid,
    input logic                              i_m_axil_arready,
    input logic [DATA_WIDTH-1:0]             i_m_axil_rdata,
    input logic [1:0]                        i_m_axil_rresp,
    input logic                              i_m_axil_rvalid,
    output logic                             i_m_axil_rready,

    output logic[ADDR_WIDTH-1:0]             d_m_axil_awaddr,
    output logic[2:0]                        d_m_axil_awprot,
    output logic                             d_m_axil_awvalid,
    input logic                              d_m_axil_awready,
    output logic[DATA_WIDTH-1:0]             d_m_axil_wdata,
    output logic[STRB_WIDTH-1:0]             d_m_axil_wstrb,
    output logic                             d_m_axil_wvalid,
    input logic                              d_m_axil_wready,
    input logic [1:0]                        d_m_axil_bresp,
    input logic                              d_m_axil_bvalid,
    output logic                             d_m_axil_bready,
    output logic[ADDR_WIDTH-1:0]             d_m_axil_araddr,
    output logic[2:0]                        d_m_axil_arprot,
    output logic                             d_m_axil_arvalid,
    input logic                              d_m_axil_arready,
    input logic [DATA_WIDTH-1:0]             d_m_axil_rdata,
    input logic [1:0]                        d_m_axil_rresp,
    input logic                              d_m_axil_rvalid,
    output logic                             d_m_axil_rready
);

axi_axil_adapter IAdapter 
(
    .clk(),
    .rst(),
    .
    .s_axi_awid(),
    .s_axi_awaddr(),
    .s_axi_awlen(),
    .s_axi_awsize(),
    .s_axi_awburst(),
    .s_axi_awlock(),
    .s_axi_awcache(),
    .s_axi_awprot(),
    .s_axi_awvalid(),
    .s_axi_awready(),
    .s_axi_wdata(),
    .s_axi_wstrb(),
    .s_axi_wlast(),
    .s_axi_wvalid(),
    .s_axi_wready(),
    .s_axi_bid(),
    .s_axi_bresp(),
    .s_axi_bvalid(),
    .s_axi_bready(),
    .s_axi_arid(),
    .s_axi_araddr(),
    .s_axi_arlen(),
    .s_axi_arsize(),
    .s_axi_arburst(),
    .s_axi_arlock(),
    .s_axi_arcache(),
    .s_axi_arprot(),
    .s_axi_arvalid(),
    .s_axi_arready(),
    .s_axi_rid(),
    .s_axi_rdata(),
    .s_axi_rresp(),
    .s_axi_rlast(),
    .s_axi_rvalid(),
    .s_axi_rready(),
    .
    .m_axil_awaddr(),
    .m_axil_awprot(),
    .m_axil_awvalid(),
    .m_axil_awready(),
    .m_axil_wdata(),
    .m_axil_wstrb(),
    .m_axil_wvalid(),
    .m_axil_wready(),
    .m_axil_bresp(),
    .m_axil_bvalid(),
    .m_axil_bready(),
    .m_axil_araddr(),
    .m_axil_arprot(),
    .m_axil_arvalid(),
    .m_axil_arready(),
    .m_axil_rdata(),
    .m_axil_rresp(),
    .m_axil_rvalid(),
    .m_axil_rready()
);

VexRiscvAxi4 #(
    .PROGADDR_RESET(32'h0201_0000)
) VexCPU (
    .timerInterrupt(?),
    .externalInterrupt(?),
    .softwareInterrupt(?),
    .debug_bus_cmd_valid(?),
    .debug_bus_cmd_ready(?),
    .debug_bus_cmd_payload_wr(?),
    .debug_bus_cmd_payload_address(?),
    .debug_bus_cmd_payload_data(?),
    .debug_bus_rsp_data(?),
    .debug_resetOut(?),
    
    .iBusAxi_ar_valid(),
    .iBusAxi_ar_ready(),
    .iBusAxi_ar_payload_addr(),
    .iBusAxi_ar_payload_id(),
    .iBusAxi_ar_payload_region(),
    .iBusAxi_ar_payload_len(),
    .iBusAxi_ar_payload_size(),
    .iBusAxi_ar_payload_burst(),
    .iBusAxi_ar_payload_lock(),
    .iBusAxi_ar_payload_cache(),
    .iBusAxi_ar_payload_qos(),
    .iBusAxi_ar_payload_prot(),
    .iBusAxi_r_valid(),
    .iBusAxi_r_ready(),
    .iBusAxi_r_payload_data(),
    .iBusAxi_r_payload_id(),
    .iBusAxi_r_payload_resp(),
    .iBusAxi_r_payload_last(),
    .dBusAxi_aw_valid(),
    .dBusAxi_aw_ready(),
    .dBusAxi_aw_payload_addr(),
    .dBusAxi_aw_payload_id(),
    .dBusAxi_aw_payload_region(),
    .dBusAxi_aw_payload_len(),
    .dBusAxi_aw_payload_size(),
    .dBusAxi_aw_payload_burst(),
    .dBusAxi_aw_payload_lock(),
    .dBusAxi_aw_payload_cache(),
    .dBusAxi_aw_payload_qos(),
    .dBusAxi_aw_payload_prot(),
    .dBusAxi_w_valid(),
    .dBusAxi_w_ready(),
    .dBusAxi_w_payload_data(),
    .dBusAxi_w_payload_strb(),
    .dBusAxi_w_payload_last(),
    .dBusAxi_b_valid(),
    .dBusAxi_b_ready(),
    .dBusAxi_b_payload_id(),
    .dBusAxi_b_payload_resp(),
    .dBusAxi_ar_valid(),
    .dBusAxi_ar_ready(),
    .dBusAxi_ar_payload_addr(),
    .dBusAxi_ar_payload_id(),
    .dBusAxi_ar_payload_region(),
    .dBusAxi_ar_payload_len(),
    .dBusAxi_ar_payload_size(),
    .dBusAxi_ar_payload_burst(),
    .dBusAxi_ar_payload_lock(),
    .dBusAxi_ar_payload_cache(),
    .dBusAxi_ar_payload_qos(),
    .dBusAxi_ar_payload_prot(),
    .dBusAxi_r_valid(),
    .dBusAxi_r_ready(),
    .dBusAxi_r_payload_data(),
    .dBusAxi_r_payload_id(),
    .dBusAxi_r_payload_resp(),
    .dBusAxi_r_payload_last(),
    .clk(),
    .reset(),
    .debugReset()
);
    
endmodule