module Channel (
    
);
    
endmodule